library verilog;
use verilog.vl_types.all;
entity ControleSemaforo_vlg_sample_tst is
    port(
        clear           : in     vl_logic;
        clock           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end ControleSemaforo_vlg_sample_tst;
