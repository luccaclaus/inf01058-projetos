library verilog;
use verilog.vl_types.all;
entity ControleSemaforo_vlg_vec_tst is
end ControleSemaforo_vlg_vec_tst;
