library verilog;
use verilog.vl_types.all;
entity Neander is
    port(
        CARGA_REM       : out    vl_logic;
        CARGA_RI        : out    vl_logic;
        clock_in        : in     vl_logic;
        clear           : in     vl_logic;
        step_button     : in     vl_logic;
        step_mode_switch: in     vl_logic;
        READ            : out    vl_logic;
        SEL             : out    vl_logic;
        PC_OUT          : out    vl_logic_vector(7 downto 0);
        INCREMENTA_PC   : out    vl_logic;
        CARGA_PC        : out    vl_logic;
        flag_N          : out    vl_logic;
        ULA_ADD         : out    vl_logic;
        ULA_AND         : out    vl_logic;
        ULA_OR          : out    vl_logic;
        ULA_NOT         : out    vl_logic;
        ULA_Y           : out    vl_logic;
        AC_OUT          : out    vl_logic_vector(7 downto 0);
        CARGA_AC        : out    vl_logic;
        CARGA_NZ        : out    vl_logic;
        flag_Z          : out    vl_logic;
        HLT             : out    vl_logic;
        GOTO_t0         : out    vl_logic;
        WRITE           : out    vl_logic;
        CARGA_RDM       : out    vl_logic;
        PC_A0           : out    vl_logic;
        PC_B0           : out    vl_logic;
        PC_C0           : out    vl_logic;
        PC_D0           : out    vl_logic;
        PC_E0           : out    vl_logic;
        PC_F0           : out    vl_logic;
        PC_G0           : out    vl_logic;
        PC_A1           : out    vl_logic;
        PC_B1           : out    vl_logic;
        PC_C1           : out    vl_logic;
        PC_D1           : out    vl_logic;
        PC_E1           : out    vl_logic;
        PC_F1           : out    vl_logic;
        PC_G1           : out    vl_logic;
        AC_A0           : out    vl_logic;
        AC_B0           : out    vl_logic;
        AC_C0           : out    vl_logic;
        AC_D0           : out    vl_logic;
        AC_E0           : out    vl_logic;
        AC_F0           : out    vl_logic;
        AC_G0           : out    vl_logic;
        AC_A1           : out    vl_logic;
        AC_B1           : out    vl_logic;
        AC_C1           : out    vl_logic;
        AC_D1           : out    vl_logic;
        AC_E1           : out    vl_logic;
        AC_F1           : out    vl_logic;
        AC_G1           : out    vl_logic
    );
end Neander;
